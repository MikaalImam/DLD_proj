`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/27/2024 04:56:47 PM
// Design Name: 
// Module Name: sprite
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// This module displays a 64x64 sprite (a dino) at the specified location on the screen
//
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module sprite_display (
    input wire clk,
    input wire reset,
    input [9:0] x_desired, y_desired,  // Position where the sprite should be displayed
    input [9:0] x, y,                   // Current x, y pixel coordinates
    output [13:0] spriteData,           // Pixel color data (RGB)
    output display_sprite               // Whether to display the sprite at the location
);

    // Define a 64x64 sprite (bicycle)
    //reg [31:0] sprite[31:0]; 
    reg [63:0] sprite[63:0];// A 64x64 sprite, 64 rows of 64 bits each
    
    initial begin
        // Define the sprite pattern for the dino
    sprite[0] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[1] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[2] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[3] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[4] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[5] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[6] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[7] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[8] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[9] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[10] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[11] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[12] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[13] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[14] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[15] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[16] = 64'b0000000000000011111111111100000000000000000000000000000000000000;
    sprite[17] = 64'b0000000000000011111111111100000000000000000000000000000000000000;
    sprite[18] = 64'b0000000000000011000000001100000000000000110011000000000000000000;
    sprite[19] = 64'b0000000000000011000000001100000000000000110011000000000000000000;
    sprite[20] = 64'b0000000000000000110000111100000000000000001111000000000000000000;
    sprite[21] = 64'b0000000000000000110000111100000000000000001111000000000000000000;
    sprite[22] = 64'b0000000000000000000000111111111111111111111100000000000000000000;
    sprite[23] = 64'b0000000000000000000000111111111111111111111100000000000000000000;
    sprite[24] = 64'b0000000000000000000011111100000000000000111111000000000000000000;
    sprite[25] = 64'b0000000000000000000011111100000000000000111111000000000000000000;
    sprite[26] = 64'b0000000000000000000011001100000000000000110011000000000000000000;
    sprite[27] = 64'b0000000000000000000011001100000000000000110011000000000000000000;
    sprite[28] = 64'b0000000000111111111111000011000000000011110011111111110000000000;
    sprite[29] = 64'b0000000000111111111111000011000000000011110011111111110000000000;
    sprite[30] = 64'b0000000011000000000011000011110000000000001100000000001100000000;
    sprite[31] = 64'b0000000011000000000011000011110000000000001100000000001100000000;
    sprite[32] = 64'b0000001111000000000011110000110000001100111100000000001111000000;
    sprite[33] = 64'b0000001111000000000011110000110000001100111100000000001111000000;
    sprite[34] = 64'b0000111100000000000000111100111100111111110000000000000011110000;
    sprite[35] = 64'b0000111100000000000000111100111100111111110000000000000011110000;
    sprite[36] = 64'b0000110000000000000000001100000011110011000000000000000000110000;
    sprite[37] = 64'b0000110000000000000000001100000011110011000000000000000000110000;
    sprite[38] = 64'b0000110000000000000000001100000011111111000000000000000000110000;
    sprite[39] = 64'b0000110000000000000000001100000011111111000000000000000000110000;
    sprite[40] = 64'b0000001100000000000000110000000000000000110000000000000011000000;
    sprite[41] = 64'b0000001100000000000000110000000000000000110000000000000011000000;
    sprite[42] = 64'b0000001111000000000011110000000000000000111100000000001111000000;
    sprite[43] = 64'b0000001111000000000011110000000000000000111100000000001111000000;
    sprite[44] = 64'b0000000011000000000011000000000000000000001100000000001100000000;
    sprite[45] = 64'b0000000011000000000011000000000000000000001100000000001100000000;
    sprite[46] = 64'b0000000000111111111100000000000000000000000011111111110000000000;
    sprite[47] = 64'b0000000000111111111100000000000000000000000011111111110000000000;
    sprite[48] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[49] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[50] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[51] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[52] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[53] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[54] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[55] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[56] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[57] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[58] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[59] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[60] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[61] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[62] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    sprite[63] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
end
        

   // Vertical positioning: map y to a sprite row
    //wire [4:0] spriteRow;
    wire [5:0] spriteRow;
    assign spriteRow = y - y_desired;  // Relative y position within the sprite, should be between 0 and 15
    // Horizontal positioning: map x to a column within the sprite row
    //wire [4:0] spriteCol;
    wire [5:0] spriteCol;
    assign spriteCol = x - x_desired;  // Relative x position within the sprite row, should be between 0 and 15
    // Get the pixel value from the sprite
    assign spriteData = (sprite[spriteRow][spriteCol] == 1'b1) ? 12'hFFF : 12'h000;  // If pixel is on, set to white; else black


    // Output the pixel value based on x, y coordinates
    assign horizontalOn = (x >= x_desired && x < x_desired + 10'd64) ? 1 : 0; //Assert horizontalOn for 7 more pixels from desired X
    assign verticalOn = (y >= y_desired && y < y_desired + 10'd64) ? 1 : 0; //Assert verticalOn for 15 more pixels from desired Y
    assign display_sprite = horizontalOn && verticalOn; //content of ROM should be displayed at these desired X,Y range
endmodule
